// ----------------------------------------------------------------------------
//
// Multi-Dataflow Composer tool - Platform Composer
// Counter module 
// Date: 2014/04/30 12:15:58
//
// ----------------------------------------------------------------------------

// ----------------------------------------------------------------------------
// Module Interface
// ----------------------------------------------------------------------------
module Cnt(
	clk,		// system clock
	reset,		// system reset
	clear,		// clear count
	maxValue,	// maximum count
	go,		// enable count
	endcount,	// finish count
	count		// count value
);
// ----------------------------------------------------------------------------

// ----------------------------------------------------------------------------
// Module Parameter(s)
// ----------------------------------------------------------------------------
parameter SIZECOUNT = 5;
// ----------------------------------------------------------------------------

// ----------------------------------------------------------------------------
// Module Signals
// ----------------------------------------------------------------------------
// Input(s)
input 				clk; 
input				reset;
input 				go;
input				clear;
input [SIZECOUNT-1 : 0]		maxValue;
// Output(s)
output [SIZECOUNT-1 : 0]	count;
output 				endcount;
// Wire(s) and Reg(s)
wire  				clk;
wire				reset;
wire 				go;
wire				clear;
wire [SIZECOUNT-1 : 0]		maxValue;
reg [SIZECOUNT-1 : 0] 		count;
reg endcount;
// ----------------------------------------------------------------------------

// ----------------------------------------------------------------------------
// Body
// ----------------------------------------------------------------------------
// Count Update
always @ (posedge clk or posedge reset)
	if (reset) 
		count <= 0;
	else if (clear)
		count <= 0;
	else if (count==maxValue)
		count <= count;
	else if (go)
		count <= count+1;

// Finish Count
always @ (count, maxValue)
	if (count==maxValue) 
		endcount <= 1;
	else 
		endcount <= 0;
// ----------------------------------------------------------------------------
		
endmodule		
// ----------------------------------------------------------------------------
// ----------------------------------------------------------------------------
// ----------------------------------------------------------------------------
