// ----------------------------------------------------------------------------
//
// Multi-Dataflow Composer tool - Platform Composer
// Register module 
// Date: 2014/04/30 12:15:58
//
// ----------------------------------------------------------------------------

// ----------------------------------------------------------------------------
// Module Interface
// ----------------------------------------------------------------------------
module Reg (
	clk,			// system clock
	enable,			// enable
	reset,			// system reset
	clear, 			// internal clear
	datain,			// input data
	dataout			// output data
);
// ----------------------------------------------------------------------------

// ----------------------------------------------------------------------------
// Module Parameter(s)
// ----------------------------------------------------------------------------
parameter SIZEDATA = 32;
// ----------------------------------------------------------------------------

// ----------------------------------------------------------------------------
// Module Signals
// ----------------------------------------------------------------------------
// Input(s)
input 			clk;
input			reset;
input 			enable;
input			clear;
input [SIZEDATA-1 : 0]	datain;
// Output(s)
output [SIZEDATA-1 : 0] dataout;
// Wire(s) and Reg(s)
wire  			clk;
wire			reset;
wire 			enable;
wire			clear;
wire [SIZEDATA-1 : 0] 	datain;
reg [SIZEDATA-1 : 0] 	dataout;
// ----------------------------------------------------------------------------

// ----------------------------------------------------------------------------
// Body
// ----------------------------------------------------------------------------
// Register
always @ (posedge clk or posedge reset) begin
	if (reset) 
		dataout <= 0;
	else if (clear) 
		dataout <=0;
	else if(enable) 
		dataout <= datain;
end
// ----------------------------------------------------------------------------
		
endmodule		
// ----------------------------------------------------------------------------
// ----------------------------------------------------------------------------
// ----------------------------------------------------------------------------
